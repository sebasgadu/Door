`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:13:04 11/08/2015 
// Design Name: 
// Module Name:    i2c_controller 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
// Modulo i2c para escribir los datos en la SDA hacia 
//////////////////////////////////////////////////////////////////////////////////
module i2c_controllerN(
       input  clk,
       inout i2c_sclk,
       inout  i2c_sdat,
       input  start,
       input reset,
       output done
    );

//Direción del SRF02 para escribir
parameter reg[7:0] address = 8'hE0;
//write de la dirección del command register
parameter reg[7:0] command_register = 8'b0;
//command que se le escribe al command register
parameter reg[7:0] command = 8'h51;
//parameter reg [23:0] i2c_data = {address,command_register, command};
parameter reg [23:0] data={address,command_register, command};

reg resetflag=1'b0;


reg [4:0] stage;
reg [6:0] sclk_divider;
reg clock_en = 1'b0;

// don't toggle the clock unless we're sending data
// clock will also be kept high when sending START and STOP symbols
assign i2c_sclk = (!clock_en) || sclk_divider[6];
wire midlow = (sclk_divider == 7'h1f);

reg sdat = 1'b1;
// rely on pull-up resistor to set SDAT high
assign i2c_sdat = (sdat) ? 1'bz : 1'b0;

reg [2:0] acks;

parameter LAST_STAGE = 5'd29;

assign ack = (acks == 3'b000);
assign done = (stage == LAST_STAGE)&&(!resetflag);


		
	
always @(posedge clk) begin
	if (reset) begin
		  sclk_divider <= 7'd0;
        stage <= LAST_STAGE;
        clock_en <= 1'b0;
        sdat <= 1'b1;
		  resetflag<=1'b1;
	end
    if (start) begin
        sclk_divider <= 7'd0;
        stage <= 5'd0;
        clock_en <= 1'b0;
        sdat <= 1'b1;
        acks <= 3'b111;
        //data <= i2c_data;
	     resetflag<=1'b0;
    end else begin
        if (sclk_divider == 7'd127) begin
            sclk_divider <= 7'd0;
            if (stage != LAST_STAGE)begin
                stage <= stage + 1'b1;
				end else resetflag <= 1'b1;

            case (stage)
                // after start
                5'd0:  clock_en <= 1'b1;
                // receive acks
                5'd9:  acks[0] <= i2c_sdat;
                5'd18: acks[1] <= i2c_sdat;
                5'd27: acks[2] <= i2c_sdat;
                // before stop
                5'd28: clock_en <= 1'b0;
            endcase
        end else
            sclk_divider <= sclk_divider + 1'b1;

        if (midlow) begin
            case (stage)
                // start
                5'd0:  sdat <= 1'b0;
                // byte 1
                5'd1:  sdat <= data[23];
                5'd2:  sdat <= data[22];
                5'd3:  sdat <= data[21];
                5'd4:  sdat <= data[20];
                5'd5:  sdat <= data[19];
                5'd6:  sdat <= data[18];
                5'd7:  sdat <= data[17];
                5'd8:  sdat <= data[16];
                // ack 1
                5'd9:  sdat <= 1'b1;
                // byte 2
                5'd10: sdat <= data[15];
                5'd11: sdat <= data[14];
                5'd12: sdat <= data[13];
                5'd13: sdat <= data[12];
                5'd14: sdat <= data[11];
                5'd15: sdat <= data[10];
                5'd16: sdat <= data[9];
                5'd17: sdat <= data[8];
                // ack 2
                5'd18: sdat <= 1'b1;
                // byte 3
                5'd19: sdat <= data[7];
                5'd20: sdat <= data[6];
                5'd21: sdat <= data[5];
                5'd22: sdat <= data[4];
                5'd23: sdat <= data[3];
                5'd24: sdat <= data[2];
                5'd25: sdat <= data[1];
                5'd26: sdat <= data[0];
                // ack 3
                5'd27: sdat <= 1'b1;
                // stop
                5'd28: sdat <= 1'b0;
                5'd29: sdat <= 1'b1;								
            endcase
        end
    end

end

endmodule

